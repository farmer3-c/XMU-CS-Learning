module binbcd4(
    input wire [3:0] b,
    output wire [4:0] p
);
    // 十位高位 (BCD码十位的最高位) - 当数值≥10时置1
    assign p[4] = (b[3] & b[2] )| (b[3] & ~b[2]&b[1]);  // b >= 10 (1010~1111)
    
    // 十位低位 (BCD码十位的最低位) - 当数值为8或9时置1
    assign p[3] = b[3] & ~b[2]&~b[1];  // 1000或1001
    
    // 个位高位 (BCD码个位的最高位)
    assign p[2] =  ( ~ b[3] & b[2]) | (b[3] & b[2] & b[1]);        // 12,14: 取0
    
    // 个位中间位
    assign p[1] = (~b[3] & b[1]) |              // 0-7: 直接取b[1]
                  (b[3] & b[2] & ~b[1]) ;        // 10,11: 置1
    
    // 个位最低位 (直接等于输入最低位)
    assign p[0] = b[0];
endmodule
